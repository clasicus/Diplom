library verilog;
use verilog.vl_types.all;
entity pwm_ver_vlg_tst is
end pwm_ver_vlg_tst;
