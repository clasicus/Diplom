library verilog;
use verilog.vl_types.all;
entity SYS_REST_vlg_tst is
end SYS_REST_vlg_tst;
