library verilog;
use verilog.vl_types.all;
entity AD7687_vlg_tst is
end AD7687_vlg_tst;
